module down_from_9 (
    output [4:0] count,

    input [3:0] set,
    input [3:0] reset,

    input clock
);


endmodule