//! Decodes binary code to output display
//!
//! See:
//!     ``display.md`` for more information.
//!
module display_decoder(
    output a, output b, output c,
    output d, output e, output f,
    output g,

    input [3:0] data
);


endmodule
