module down_from_5 (
    output [3:0] count,

    input [2:0] set,
    input [2:0] reset,

    input clock
);


endmodule